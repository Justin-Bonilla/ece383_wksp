------
-- Lt Col James Trimble, 15 Jan 2025
-- Generates VGA signal with graphics
------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.ece383_pkg.ALL;
 
entity vga is
	Port(	clk: in  STD_LOGIC;
			reset_n : in  STD_LOGIC;
			vga : out vga_t;
            pixel : out pixel_t;
			trigger : in trigger_t;
            ch1 : in channel_t;
            ch2 : in channel_t);
end vga;

architecture vga_arch of vga is
		signal current_pos : coordinate_t;
		
	
begin

vga_sig_gen : vga_signal_generator
port map(
    clk      => clk,
    reset_n  => reset_n,
    position => current_pos,
    vga      => vga
);

pixel.coordinate <= current_pos;
--pixel_position <= current_pos;

col_map : color_mapper
port map(  color => pixel.color,
           position => current_pos, --pixel_position,
		   trigger => trigger,
           ch1 => ch1,
           ch2 => ch2
);

end vga_arch;
